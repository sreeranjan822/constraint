class







endclass
