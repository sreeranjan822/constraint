class

function





endclass
